library ieee;
use ieee.std_logic_1164.all;
library work;
use work.Gates.all;

entity one2eight  is
  port (d: in std_logic_vector(15 downto 0);s: in std_logic_vector(2 downto 0); y0: out std_logic_vector(15 downto 0); y1: out std_logic_vector(15 downto 0); y2: out std_logic_vector(15 downto 0); y3: out std_logic_vector(15 downto 0); y4: out std_logic_vector(15 downto 0); y5: out std_logic_vector(15 downto 0); y6: out std_logic_vector(15 downto 0); y7: out std_logic_vector(15 downto 0));
end entity one2eight;

architecture Struct of one2eight is

begin
    y0 <= (((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))&((not s(0)) and (not s(1)) and (not s(2)))) and d;
    y1 <= (((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))&((s(0)) and (not s(1)) and (not s(2)))) and d;
    y2 <= (((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))&((not s(0)) and (s(1)) and (not s(2)))) and d;
    y3 <= (((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))&((s(0)) and (s(1)) and (not s(2)))) and d;
    y4 <= (((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))&((not s(0)) and (not s(1)) and (s(2)))) and d;
    y5 <= (((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))&((s(0)) and (not s(1)) and (s(2)))) and d;
    y6 <= (((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))&((not s(0)) and (s(1)) and (s(2)))) and d;
    y7 <= (((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))&((s(0)) and (s(1)) and (s(2)))) and d;

end Struct;